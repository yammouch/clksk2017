module stimulus (
 input             RSTX,
 input             CLK,
 input             RSTXF,
 input             CLKF,
 input             CLKF_DATA,
 input             RSTXS,
 input             CLKS,
 input             CLKSS,
 input             CLR,
 input             SERDESSTROBE,
 input      [ 7:0] MAIN_MODE,
 input      [ 7:0] SUB_MODE,
 output reg [30:0] CTRL,
 output     [ 1:0] DOUT,
 input      [ 1:0] DIN,
 output            PHY_INIT,
 output     [59:0] RECV_CNT,
 output     [63:0] ERR_CNT);

always @(posedge CLK)
  case (MAIN_MODE)
  8'd1 : DOUT <= 30'b1111_01_0000_00_0000_00_0000_0000_1000;
  8'd2 : DOUT <= 30'b1111_01_0000_00_0000_00_0000_0000_0000;
  8'd3 : DOUT <= 30'b1111_10_0000_00_0000_00_0000_0000_0010;
  8'd4 : DOUT <= 30'b1111_10_0000_00_0000_00_0000_0000_0000;
  8'd5 : begin
    DOUT[29:26] <= 4'b1111;
    DOUT[   25] <= SUB_MODE[0];
    DOUT[24: 0] <= 25'b1_0000_00_0000_00_0000_0000_0000;
  end
  8'd6 : begin
    DOUT[29:25] <= 5'b1111_1;
    DOUT[   25] <= SUB_MODE[0];
    DOUT[24: 0] <= 24'b0000_00_0000_00_0000_0000_0000;
  end
  8'd7 : begin
    DOUT[29:20] <= 10'b0000_00_1111;
    DOUT[19:18] <= {2{SUB_MODE[0]}};
    DOUT[17: 0] <= 18'b0000_00_0000_0000_0000;
  end
  8'd8 : DOUT <= 30'b0000_00_1111_11_0000_00_0000_0000_0000;
  8'd9 : DOUT <= 30'b0000_00_1111_11_0000_00_0000_0000_0000;
  8'd10: DOUT <= 30'b0111_01_0000_11_0000_00_0000_0000_0000;
  8'd11: DOUT <= 30'b0111_01_0000_11_0000_00_0000_0000_0000;
  8'd12: DOUT <= 30'b0111_01_0000_11_0000_00_0000_0000_0000;
  8'd13: DOUT <= 30'b0000_00_0000_11_0000_00_0000_0000_0000;
  8'd14: DOUT <= 30'b0000_00_0100_11_0000_00_0000_0000_0000;
  8'd15: DOUT <= 30'b0000_00_1000_11_0000_00_0000_0000_0000;
  8'd16: DOUT <= 30'b0000_00_1100_11_0000_00_0000_0000_0000;
  8'd17: DOUT <= 30'b0000_00_0000_11_0000_00_0000_0000_0000;
  8'd18: DOUT <= 30'b0000_00_0001_11_0000_00_0000_0000_0000;
  8'd19: DOUT <= 30'b0000_00_0010_11_0000_00_0000_0000_0000;
  8'd20: DOUT <= 30'b0000_00_0011_11_0000_00_0000_0000_0000;
  8'd21: DOUT <= 30'b0101_01_1100_10_0000_00_0000_0000_0000;
  8'd22: DOUT <= 30'b1010_10_0011_01_0000_00_0000_0000_0000;
  8'd23: DOUT <= 30'b0101_01_0000_10_0000_00_0000_0000_0000;
  8'd24: DOUT <= 30'b0101_01_0100_10_0000_00_0000_0000_0000;
  8'd25: DOUT <= 30'b0101_01_1000_10_0000_00_0000_0000_0000;
  8'd26: DOUT <= 30'b0101_01_1100_10_0000_00_0000_0000_0000;
  8'd27: DOUT <= 30'b1010_10_0000_01_0000_00_0000_0000_0000;
  8'd28: DOUT <= 30'b1010_10_0001_01_0000_00_0000_0000_0000;
  8'd29: DOUT <= 30'b1010_10_0010_01_0000_00_0000_0000_0000;
  8'd30: DOUT <= 30'b1010_10_0011_01_0000_00_0000_0000_0000;
  8'd31: DOUT <= 30'b0000_00_1111_11_0000_00_0000_0000_0000;
  8'd32: DOUT <= 30'b1111_00_0000_00_0000_00_0000_0000_0000;
  8'd33: DOUT <= 30'b1111_00_0000_00_0100_00_0000_0000_0000;
  8'd34: DOUT <= 30'b1111_00_0000_00_1000_00_0000_0000_0000;
  8'd35: DOUT <= 30'b1111_00_0000_00_1100_00_0000_0000_0000;
  8'd36: DOUT <= 30'b1111_00_0000_00_0100_10_0000_0000_0000;
  8'd37: DOUT <= 30'b1111_00_0000_00_1000_10_0000_0000_0000;
  8'd38: DOUT <= 30'b1111_00_0000_00_1100_10_0000_0000_0000;
  8'd39: DOUT <= 30'b1111_00_0000_00_0000_00_0000_0000_0000;
  8'd40: DOUT <= 30'b1111_00_0000_00_0001_00_0000_0000_0000;
  8'd41: DOUT <= 30'b1111_00_0000_00_0010_00_0000_0000_0000;
  8'd42: DOUT <= 30'b1111_00_0000_00_0011_00_0000_0000_0000;
  8'd43: DOUT <= 30'b1111_00_0000_00_0001_01_0000_0000_0000;
  8'd44: DOUT <= 30'b1111_00_0000_00_0010_01_0000_0000_0000;
  8'd45: DOUT <= 30'b1111_00_0000_00_0011_01_0000_0000_0000;
  8'd46: begin
    DOUT[29:6] <= 24'b1111_00_0000_00_0000_00_0010_00;
    DOUT[   5] <= SUB_MODE[0];
    DOUT[ 4:0] <= 5'b0_0000;
  end
  8'd47: begin
    DOUT[29:5] <= 25'b1111_00_0000_00_0000_00_0010_00_0;
    DOUT[   4] <= SUB_MODE[0];
    DOUT[ 3:0] <= 4'b0000;
  end
  8'd48: DOUT <= 30'b1111_00_0000_00_0000_00_0000_0000_1000;
  8'd49: DOUT <= 30'b1111_00_0000_00_0100_00_0000_0000_1000;
  8'd50: DOUT <= 30'b1111_00_0000_00_1000_00_0000_0000_1000;
  8'd51: DOUT <= 30'b1111_00_0000_00_1100_00_0000_0000_1000;
  8'd52: DOUT <= 30'b1111_00_0000_00_0100_10_0000_0000_1000;
  8'd53: DOUT <= 30'b1111_00_0000_00_1000_10_0000_0000_1000;
  8'd54: DOUT <= 30'b1111_00_0000_00_1100_10_0000_0000_1000;
  8'd55: DOUT <= 30'b1111_00_0000_00_0000_00_0000_0000_0010;
  8'd56: DOUT <= 30'b1111_00_0000_00_0001_00_0000_0000_0010;
  8'd57: DOUT <= 30'b1111_00_0000_00_0010_00_0000_0000_0010;
  8'd58: DOUT <= 30'b1111_00_0000_00_0011_00_0000_0000_0010;
  8'd59: DOUT <= 30'b1111_00_0000_00_0001_01_0000_0000_0010;
  8'd60: DOUT <= 30'b1111_00_0000_00_0010_01_0000_0000_0010;
  8'd61: DOUT <= 30'b1111_00_0000_00_0011_01_0000_0000_0010;
  8'd62: begin
    DOUT[29:8] <= 22'b1111_00_0000_00_0000_00_0010;
    DOUT[   7] <= SUB_MODE[0];
    DOUT[ 6:0] <= 7'b000_1000;
  end
  8'd63: begin
    DOUT[29:7] <= 23'b1111_00_0000_00_0000_00_0001_0;
    DOUT[   6] <= SUB_MODE[0];
    DOUT[ 5:0] <= 6'b00_0010;
  end
  endcase
  8'd64: DOUT <= 30'b1000_00_1100_00_0000_00_0000_0000_0000;
  8'd65: DOUT <= 30'b1000_00_1100_00_0000_00_0000_0000_0100;
  8'd66: DOUT <= 30'b0100_00_0011_00_0000_00_0000_0000_0000;
  8'd67: DOUT <= 30'b0100_00_0011_00_0000_00_0000_0000_0001;
  8'd68: DOUT <= 30'b0010_00_0000_10_1100_00_0000_0000_0000;
  8'd69: DOUT <= 30'b0001_00_0000_01_0011_00_0000_0000_0000;
  default: DOUT <= 30'd0;

endmodule
