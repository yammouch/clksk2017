module stimulus (
 input             RSTX,
 input             CLK,
 input             RSTXF,
 input             CLKF,
 input             CLKF_DATA,
 input             RSTXS,
 input             CLKS,
 input             CLKSS,
 input             CLR,
 input             SERDESSTROBE,
 input      [ 7:0] MAIN_MODE,
 input      [ 7:0] SUB_MODE,
 output reg [30:0] CTRL,
 output     [ 1:0] DOUT,
 input      [ 1:0] DIN,
 output            PHY_INIT,
 output     [59:0] RECV_CNT,
 output     [63:0] ERR_CNT);

assign RECV_CNT = 60'd0;
assign ERR_CNT  = 64'd0;
assign PHY_INIT = 1'b0;

always @(posedge CLKF) CTRL[0] <= 1'b0;

always @(posedge CLKF)
  case (MAIN_MODE)
  8'd1 : CTRL[30:1] <= 30'b1111_01_0000_00_0000_00_0000_0000_1000;
  8'd2 : CTRL[30:1] <= 30'b1111_01_0000_00_0000_00_0000_0000_0000;
  8'd3 : CTRL[30:1] <= 30'b1111_10_0000_00_0000_00_0000_0000_0010;
  8'd4 : CTRL[30:1] <= 30'b1111_10_0000_00_0000_00_0000_0000_0000;
  8'd5 : begin
    CTRL[30:27] <= 4'b1111;
    CTRL[   26] <= SUB_MODE[0];
    CTRL[25: 1] <= 25'b1_0000_00_0000_00_0000_0000_0000;
  end
  8'd6 : begin
    CTRL[30:27] <= 5'b1111_1;
    CTRL[   26] <= SUB_MODE[0];
    CTRL[25: 1] <= 24'b0000_00_0000_00_0000_0000_0000;
  end
  8'd7 : begin
    CTRL[30:21] <= 10'b0000_00_1111;
    CTRL[20:19] <= {2{SUB_MODE[0]}};
    CTRL[18: 1] <= 18'b0000_00_0000_0000_0000;
  end
  8'd8 : CTRL[30:1] <= 30'b0000_00_1111_11_0000_00_0000_0000_0000;
  8'd9 : CTRL[30:1] <= 30'b0000_00_1111_11_0000_00_0000_0000_0000;
  8'd10: CTRL[30:1] <= 30'b0111_01_0000_11_0000_00_0000_0000_0000;
  8'd11: CTRL[30:1] <= 30'b0111_01_0000_11_0000_00_0000_0000_0000;
  8'd12: CTRL[30:1] <= 30'b0111_01_0000_11_0000_00_0000_0000_0000;
  8'd13: CTRL[30:1] <= 30'b0000_00_0000_11_0000_00_0000_0000_0000;
  8'd14: CTRL[30:1] <= 30'b0000_00_0100_11_0000_00_0000_0000_0000;
  8'd15: CTRL[30:1] <= 30'b0000_00_1000_11_0000_00_0000_0000_0000;
  8'd16: CTRL[30:1] <= 30'b0000_00_1100_11_0000_00_0000_0000_0000;
  8'd17: CTRL[30:1] <= 30'b0000_00_0000_11_0000_00_0000_0000_0000;
  8'd18: CTRL[30:1] <= 30'b0000_00_0001_11_0000_00_0000_0000_0000;
  8'd19: CTRL[30:1] <= 30'b0000_00_0010_11_0000_00_0000_0000_0000;
  8'd20: CTRL[30:1] <= 30'b0000_00_0011_11_0000_00_0000_0000_0000;
  8'd21: CTRL[30:1] <= 30'b0101_01_1100_10_0000_00_0000_0000_0000;
  8'd22: CTRL[30:1] <= 30'b1010_10_0011_01_0000_00_0000_0000_0000;
  8'd23: CTRL[30:1] <= 30'b0101_01_0000_10_0000_00_0000_0000_0000;
  8'd24: CTRL[30:1] <= 30'b0101_01_0100_10_0000_00_0000_0000_0000;
  8'd25: CTRL[30:1] <= 30'b0101_01_1000_10_0000_00_0000_0000_0000;
  8'd26: CTRL[30:1] <= 30'b0101_01_1100_10_0000_00_0000_0000_0000;
  8'd27: CTRL[30:1] <= 30'b1010_10_0000_01_0000_00_0000_0000_0000;
  8'd28: CTRL[30:1] <= 30'b1010_10_0001_01_0000_00_0000_0000_0000;
  8'd29: CTRL[30:1] <= 30'b1010_10_0010_01_0000_00_0000_0000_0000;
  8'd30: CTRL[30:1] <= 30'b1010_10_0011_01_0000_00_0000_0000_0000;
  8'd31: CTRL[30:1] <= 30'b0000_00_1111_11_0000_00_0000_0000_0000;
  8'd32: CTRL[30:1] <= 30'b1111_00_0000_00_0000_00_0000_0000_0000;
  8'd33: CTRL[30:1] <= 30'b1111_00_0000_00_0100_00_0000_0000_0000;
  8'd34: CTRL[30:1] <= 30'b1111_00_0000_00_1000_00_0000_0000_0000;
  8'd35: CTRL[30:1] <= 30'b1111_00_0000_00_1100_00_0000_0000_0000;
  8'd36: CTRL[30:1] <= 30'b1111_00_0000_00_0100_10_0000_0000_0000;
  8'd37: CTRL[30:1] <= 30'b1111_00_0000_00_1000_10_0000_0000_0000;
  8'd38: CTRL[30:1] <= 30'b1111_00_0000_00_1100_10_0000_0000_0000;
  8'd39: CTRL[30:1] <= 30'b1111_00_0000_00_0000_00_0000_0000_0000;
  8'd40: CTRL[30:1] <= 30'b1111_00_0000_00_0001_00_0000_0000_0000;
  8'd41: CTRL[30:1] <= 30'b1111_00_0000_00_0010_00_0000_0000_0000;
  8'd42: CTRL[30:1] <= 30'b1111_00_0000_00_0011_00_0000_0000_0000;
  8'd43: CTRL[30:1] <= 30'b1111_00_0000_00_0001_01_0000_0000_0000;
  8'd44: CTRL[30:1] <= 30'b1111_00_0000_00_0010_01_0000_0000_0000;
  8'd45: CTRL[30:1] <= 30'b1111_00_0000_00_0011_01_0000_0000_0000;
  8'd46: begin
    CTRL[30:7] <= 24'b1111_00_0000_00_0000_00_0010_00;
    CTRL[   6] <= SUB_MODE[0];
    CTRL[ 5:1] <= 5'b0_0000;
  end
  8'd47: begin
    CTRL[30:6] <= 25'b1111_00_0000_00_0000_00_0010_00_0;
    CTRL[   5] <= SUB_MODE[0];
    CTRL[ 4:1] <= 4'b0000;
  end
  8'd48: CTRL[30:1] <= 30'b1111_00_0000_00_0000_00_0000_0000_1000;
  8'd49: CTRL[30:1] <= 30'b1111_00_0000_00_0100_00_0000_0000_1000;
  8'd50: CTRL[30:1] <= 30'b1111_00_0000_00_1000_00_0000_0000_1000;
  8'd51: CTRL[30:1] <= 30'b1111_00_0000_00_1100_00_0000_0000_1000;
  8'd52: CTRL[30:1] <= 30'b1111_00_0000_00_0100_10_0000_0000_1000;
  8'd53: CTRL[30:1] <= 30'b1111_00_0000_00_1000_10_0000_0000_1000;
  8'd54: CTRL[30:1] <= 30'b1111_00_0000_00_1100_10_0000_0000_1000;
  8'd55: CTRL[30:1] <= 30'b1111_00_0000_00_0000_00_0000_0000_0010;
  8'd56: CTRL[30:1] <= 30'b1111_00_0000_00_0001_00_0000_0000_0010;
  8'd57: CTRL[30:1] <= 30'b1111_00_0000_00_0010_00_0000_0000_0010;
  8'd58: CTRL[30:1] <= 30'b1111_00_0000_00_0011_00_0000_0000_0010;
  8'd59: CTRL[30:1] <= 30'b1111_00_0000_00_0001_01_0000_0000_0010;
  8'd60: CTRL[30:1] <= 30'b1111_00_0000_00_0010_01_0000_0000_0010;
  8'd61: CTRL[30:1] <= 30'b1111_00_0000_00_0011_01_0000_0000_0010;
  8'd62: begin
    CTRL[30:9] <= 22'b1111_00_0000_00_0000_00_0010;
    CTRL[   8] <= SUB_MODE[0];
    CTRL[ 7:1] <= 7'b000_1000;
  end
  8'd63: begin
    CTRL[30:8] <= 23'b1111_00_0000_00_0000_00_0001_0;
    CTRL[   7] <= SUB_MODE[0];
    CTRL[ 6:1] <= 6'b00_0010;
  end
  8'd64: CTRL[30:1] <= 30'b1000_00_1100_00_0000_00_0000_0000_0000;
  8'd65: CTRL[30:1] <= 30'b1000_00_1100_00_0000_00_0000_0000_0100;
  8'd66: CTRL[30:1] <= 30'b0100_00_0011_00_0000_00_0000_0000_0000;
  8'd67: CTRL[30:1] <= 30'b0100_00_0011_00_0000_00_0000_0000_0001;
  8'd68: CTRL[30:1] <= 30'b0010_00_0000_10_1100_00_0000_0000_0000;
  8'd69: CTRL[30:1] <= 30'b0001_00_0000_01_0011_00_0000_0000_0000;
  default: CTRL[30:1] <= 30'd0;
  endcase

wire [1:0] seq_32;
seq #(.BW_SEQ(3'd2), .SEQ_CNT(2'd2), .BW_SEQ_CNT(2'd2), .RV(2'd0),
 .BW_TIMEOUT(1'b1) ) i_seq_32 (
 .RSTX(RSTXF), .CLK(CLKF), .CLR(CLR), .SEQ(seq_32),
 .PTN ( { 2'b10, 1'b0
        , 2'b01, 1'b1
        , 2'b00, 1'b1 } )
);

reg [7:0] vio_ctrl;

assign DOUT[1] = vio_ctrl[7] ? vio_ctrl[6] : 1'bz;
assign DOUT[0] = vio_ctrl[5] ? vio_ctrl[4] : 1'bz;
assign DIN[1]  = vio_ctrl[3] ? vio_ctrl[2] : 1'bz;
assign DIN[0]  = vio_ctrl[1] ? vio_ctrl[0] : 1'bz;

always @(posedge CLKF or negedge RSTXF)
  case (MAIN_MODE)
  8'd1 : vio_ctrl <= 8'b10101010_00000000;
  8'd2 : vio_ctrl <= 8'b10101010_00000000;
  8'd3 : vio_ctrl <= 8'b10101010_00000000;
  8'd4 : vio_ctrl <= 8'b1010_0000;
  8'd5 : vio_ctrl <= 8'b1010_0000;
  8'd6 : vio_ctrl <= 8'b1010_0000;
  8'd7 : vio_ctrl <= { 1'b1, seq_32[1], 1'b1, seq_32[0], 4'b0000 };
  8'd8 : vio_ctrl <= 8'b00000000;
  8'd32: vio_ctrl <= { 1'b1, seq_32[1], 1'b1, seq_32[0], 4'b0000 };
  8'd33: vio_ctrl <= { 1'b1, seq_32[1], 1'b1, seq_32[0], 4'b0000 };
  8'd34: vio_ctrl <= { 1'b1, seq_32[1], 1'b1, seq_32[0], 4'b0000 };
  8'd35: vio_ctrl <= { 1'b1, seq_32[1], 1'b1, seq_32[0], 4'b0000 };
  8'd36: vio_ctrl <= { 1'b1, seq_32[1], 1'b1, seq_32[0], 4'b0000 };
  8'd37: vio_ctrl <= { 1'b1, seq_32[1], 1'b1, seq_32[0], 4'b0000 };
  8'd38: vio_ctrl <= { 1'b1, seq_32[1], 1'b1, seq_32[0], 4'b0000 };
  8'd46: vio_ctrl <= 8'b00000000;
  8'd48: vio_ctrl <= { 4'b0000, 1'b1, seq_32[1], 1'b1, seq_32[0] };
  8'd49: vio_ctrl <= { 4'b0000, 1'b1, seq_32[1], 1'b1, seq_32[0] };
  8'd50: vio_ctrl <= { 4'b0000, 1'b1, seq_32[1], 1'b1, seq_32[0] };
  8'd51: vio_ctrl <= { 4'b0000, 1'b1, seq_32[1], 1'b1, seq_32[0] };
  8'd52: vio_ctrl <= { 4'b0000, 1'b1, seq_32[1], 1'b1, seq_32[0] };
  8'd53: vio_ctrl <= { 4'b0000, 1'b1, seq_32[1], 1'b1, seq_32[0] };
  8'd54: vio_ctrl <= { 4'b0000, 1'b1, seq_32[1], 1'b1, seq_32[0] };
  8'd62: vio_ctrl <= 8'b00000000;
  default: vio_ctrl <= 8'b00000000;
  endcase

endmodule
